zifan@zifan-Dell-System-XPS-L502X.6832:1403083494